//MACROS

//Colours
`define TRANSPARENT 16'h07e7
`define BLACK 0
`define WHITE 16'hffff
`define GREY 16'h8c71

//Menu
`define MENUTRIANGLE 16'h26bb
`define LIGHTPINK 16'hf4d0
`define LIGHTYELLOW 16'hf710
`define LIGHTPURPLE 16'hde1e
`define LIGHTBLUE 16'hdf5e
`define LIGHTORANGE 16'hf54d
`define DARKPURPLE 16'h8ada
`define DARKORANGE 16'hfc80
`define DARKPINK 16'hfb6a
`define DARKBLUE 16'h3370
`define DARKGREEN 16'h2360

//Volume Bar
`define THEME1TIER1 16'h07e0
`define THEME1TIER2 16'hffe0
`define THEME1TIER3 16'hf800

`define THEME2BORDER 16'h4a69
`define THEME2TIER1 16'h8f3d
`define THEME2TIER2 16'h34b4
`define THEME2TIER3 16'h218f

//Screem Hero
`define SCREEMBG 16'hafff
`define CATHEIGHT 13
`define CATLEGWIDTH 13 
`define CATWIDTH 16
`define BLOCKWIDTH 35

//Waveform
`define PURPLE_THEME1 16'h071F
`define PURPLE_THEME1h 16'h049F
`define PURPLE_THEME2 16'h021F
`define PURPLE_THEME2h 16'h481F
`define PURPLE_THEME3 16'hC81F
`define PURPLE_THEME3h 16'hF81A
`define PURPLE_THEME4 16'hF80E
`define PURPLE_THEME4h 16'hF800

//Big Bad Wolf
`define DYING_COLOUR 16'h1a42

//Slappy Hands
`define PLAYER1COLOUR 16'h92c1
`define PLAYER2COLOUR 16'h701f


